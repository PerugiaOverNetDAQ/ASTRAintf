library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.math_real.all;

use work.basic_package.all;
use work.ASTRApackage.all;


entity ASTRA_sim is

end entity ASTRA_sim;

architecture behav of ASTRA_sim is

begin

end architecture behav;
